library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TopLevel is
    port (
        
    );
end entity TopLevel;

architecture rtl of TopLevel is
    
begin
    
    
    
end architecture rtl;